module CPU_wrapper(



);


endmodule